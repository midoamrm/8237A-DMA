module testato(leba , teba);

input leba;
output teba;

assign teba=leba;

endmodule 
